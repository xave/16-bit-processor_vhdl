LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY CU16bit IS
PORT (	CLK:  IN STD_LOGIC ; --This is the clock that controls the entire circuit.
		Reset: IN STD_LOGIC ;
		DATA: IN STD_LOGIC_VECTOR(15 DOWNTO 0) ; --aka FUNCTIONS
		Wr: OUT STD_LOGIC; --This is the Write enable for the memory. 1=write. 0=read		)
		REG_IN: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) ; --register enable
		REG_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) ; --tristate enable
		RegA_in: OUT STD_LOGIC ;
		RegG_in: OUT_STD_LOGIC ;
		RegG_out: OUT STD_LOGIC; 
		ALU_com:  OUT STD_LOGIC_VECTOR(3 DOWNTO 0) ;
		Jmp_en: OUT STD_LOGIC ; --This lets the program counter jump. --Otherwise it increments on its own.
		jmp_addr: OUT STD_LOGIC_VECTOR(15 DOWNTO 0) ;
		Done: OUT_STD_LOGIC ; -- This tells the program counter to increment when asserted.
		Ce: OUT STD_LOGIC ) ;--This lets the ram do stuff when enabled.
END ENTITY;

ARCHITECTURE Behavior OF CU16bit IS
TYPE State_type IS (HOME, LOAD, LOAD2, LOAD3, MOV, MOV2, ADD, ADD2, ADD3, ADD4, ADD5, ADD6,  SUB, SUB2, SUB3, SUB4, SUB5, SUB6, MULT, DIV, BGTE, JMP, XOR1,  XOR2, XOR3, XOR4, XOR5, XOR6) ;
SIGNAL Y_present, Y_next : State_type ;
SIGNAL data_enable : STD_LOGIC_VECTOR(1 DOWNTO 0):="00" ;
SIGNAL Reset, Clock, DATA : STD_LOGIC ; 
SIGNAL count : std_logic_vector (7 DOWNTO 0) ;







----------------------------------------------------------------
--Process A: This tells you to either move through states or 
--           reset.
BEGIN
	PROCESS (Clock, Reset)
		BEGIN
		IF Reset = '1' THEN
			y_present <= HOME; -- resets to Home state
			sCOm<= (others=>'0') ;
		ELSIF (Clock'EVENT AND Clock = '1') THEN
			y_present <= y_next ;--next state becomes the present state 
			--DATA<= DATA ;--We needed this to keep the ALU command from overwriting each tme
		END IF ;
	END PROCESS ;

----------------------------------------------------------------
----------------------------------------------------------------

--Process B: This defines how one moves through states.

PROCESS (Y_present) -- state table
BEGIN

	CASE Y_present IS

	---------HOME---------
	WHEN HOME =>
	Done<='0' ;	
		 --declare outputs--   
	IF (DATA(15 DOWNTO 12) = "0000") THEN
		Y_next <= HOME;

	ELSIF (DATA(15 DOWNTO 12) = "0001") THEN
		Y_next <= LOAD;

	ELSIF (DATA(15 DOWNTO 12) = "0010") THEN
		Y_next <= MOV;

	ELSIF (DATA(15 DOWNTO 12) = "0011") THEN
		Y_next <= ADD;

	ELSIF (DATA(15 DOWNTO 12) = "0100") THEN
		Y_next <= SUB;

	ELSIF (DATA(15 DOWNTO 12) = "0101") THEN
		Y_next <= MULT;

	ELSIF (DATA(15 DOWNTO 12) = "0110") THEN
		Y_next <= DIV;

	ELSIF (DATA(15 DOWNTO 12) = "0111") THEN
		Y_next <= XOR1;

	ELSIF (DATA(15 DOWNTO 12) = "1000") THEN
		Y_next <= JMP;

	ELSIF (DATA(15 DOWNTO 12) = "1001") THEN
		Y_next <= BGT;

	ELSIF (DATA(15 DOWNTO 12) = "1010") THEN
		Y_next <= COM;

	END IF;
------------------------------------------------------------------------------------
     ------------------------------------LOAD---------
WHEN LOAD =>
			 --declare outputs--   
Y_next <= LOAD2;
Wr<='0';--RAM is in "read mode"
CE<='1';
Jmp_en<='1';
jmp_addr<= "00000000" & DATA(7 DOWNTO 0);

 ---------LOAD2---------
WHEN LOAD2 =>
			 --declare outputs--   
Y_next <=LOAD3;
Wr<='1';--RAM is in "Write mode."
-- find REG_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<= "0000000000000001";
END IF;
---------LOAD3---------
WHEN LOAD3 =>
			 --declare outputs--   

Y_next<=HOME;
REG_IN <= (others  => '0');
CE<='0';
Done<='1';
--------------------MOV---------------------------------------------------------
WHEN MOV =>
                         --declare outputs-- 

Y_next<=MOV2;
--Reg_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--Reg IN
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_IN<="0000000000000001";
END IF;

WHEN MOV2=>
Y_next<=HOME;
Reg_IN<= (others => '0');
Reg_OUT<= (others => '0');
Done<='1';
----------------ADD-------------------------------------------------
WHEN ADD=>
Y_next<=ADD2;
--Regx_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;

RegA_in<='1';

WHEN ADD2=>
Y_next<=ADD3;
RegA_in<='0';
Reg_OUT<= (others => '0'); 

--Regy_out--- 
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--
ALU_com<= DATA(15 DOWNTO 12);

WHEN ADD3=>   --WAIT
Y_next<= ADD4;
Reg_OUT<=(others =>'0');
ALU_com<=DATA(15 DOWNTO 12);

WHEN ADD4=>

Y_next<=ADD5;
RegG_IN<='1';
RegG_OUT<='1';

WHEN ADD5=>
y_NEXT<=ADD6;
--Regx_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<= "0000000000000001";
END IF;

WHEN ADD6=>
Y_next<=HOME;
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
RegG_IN<='0';
RegG_OUT<='0';
Done<='1';






































------SUBTRACT------------------------------------------------------
WHEN SUB=>
Y_next<=SUB2;
--Regx_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;

RegA_in<='1';

WHEN SUB2=>
Y_next<=SUB3;
RegA_in<='0';
Reg_OUT<= (others => '0'); 

--Regy_out--- 
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--
ALU_com<= DATA(15 DOWNTO 12);

WHEN SUB3=>   --WAIT
Y_next<= SUB4;
Reg_OUT<=(others =>'0');
ALU_com<=DATA(15 DOWNTO 12);

WHEN SUB4=>

Y_next<=SUB5;
RegG_IN<='1';
RegG_OUT<='1';

WHEN SUB5=>
y_NEXT<=SUB6;
--Regx_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<="0000000000000001";
END IF;

WHEN SUB6=>
Y_next<=HOME;
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
RegG_IN<='0';
RegG_OUT<='0';
Done<='1';
------compare------------------------------------------------------
WHEN CMP=>
Y_next<=CMP2;
--Regx_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;

RegA_in<='1';

WHEN CMP2=>
Y_next<=CMP3;
RegA_in<='0';
Reg_OUT<= (others => '0'); 

--Regy_out--- 
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--
ALU_com<= DATA(15 DOWNTO 12);

WHEN CMP3=>   --WAIT
Y_next<= CMP4;
Reg_OUT<=(others =>'0');
ALU_com<=DATA(15 DOWNTO 12);

WHEN CMP4=>

Y_next<=CMP5;
RegG_IN<='1';
RegG_OUT<='1';

WHEN CMP5=>
y_NEXT<=CMP6;
--Regx_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<="0000000000000001";
END IF;

WHEN CMP6=>
Y_next<=HOME;
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
RegG_IN<='0';
RegG_OUT<='0';
Done<='1';
------xor------------------------------------------------------
WHEN XOR1=>
Y_next<=XOR2;
--Regx_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;

RegA_in<='1';

WHEN XOR2=>
Y_next<=XOR3;
RegA_in<='0';
Reg_OUT<= (others => '0'); 

--Regy_out--- 
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--
ALU_com<= DATA(15 DOWNTO 12);

WHEN XOR3=>   --WAIT
Y_next<= XOR4;
Reg_OUT<=(others =>'0');
ALU_com<=DATA(15 DOWNTO 12);

WHEN XOR4=>

Y_next<=XOR1;
RegG_OUT<='1';

WHEN XOR5=>
y_NEXT<=XOR6;
--Regx_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<="0000000000000001";
END IF;

WHEN XOR6=>
Y_next<=HOME;
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
RegG_IN<='0';
RegG_OUT<='0';
Done<='1';
-----------------JUMP------------------
WHEN JMP=>
Y_next<=JMP2;
Jmp_en<='1';
Jmp_addr<= DATA(11 DOWNTO 4) & "00000000";
Wr<='0';
CE<='1';

WHEN JMP2=>
Y_next<=HOME;
Jmp_en<='0';
CE<='0';
Done<='1';





---Branch if not equal----
WHEN BGT1=>
Y_next<=BGT2;
--Regx_OUT
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;

RegA_in<='1';

WHEN BGT2=>
Y_next<=BGT3;
RegA_in<='0';
Reg_OUT<= (others => '0'); 

--Regy_out--- 
IF DATA(7 DOWNTO 4)="0000" THEN 
Reg_OUT<="1000000000000000";
ELSIF DATA(7 DOWNTO 4) ="0001" THEN
Reg_OUT<="0100000000000000";
ELSIF DATA(7 DOWNTO 4) ="0010" THEN
Reg_OUT<="0010000000000000";
ELSIF DATA(7 DOWNTO 4) ="0011" THEN
Reg_OUT<="0001000000000000";
ELSIF DATA(7 DOWNTO 4) ="0100" THEN
Reg_OUT<="0000100000000000";
ELSIF DATA(7 DOWNTO 4) ="0101" THEN
Reg_OUT<="0000010000000000";
ELSIF DATA(7 DOWNTO 4) ="0110" THEN
Reg_OUT<="0000001000000000";
ELSIF DATA(7 DOWNTO 4) ="0111" THEN
Reg_OUT<="0000000100000000";
ELSIF DATA(7 DOWNTO 4) ="1000" THEN
Reg_OUT<="0000000010000000";
ELSIF DATA(7 DOWNTO 4) ="1001" THEN
Reg_OUT<="0000000001000000";
ELSIF DATA(7 DOWNTO 4) ="1010" THEN
Reg_OUT<="0000000000100000";
ELSIF DATA(7 DOWNTO 4) ="1011" THEN
Reg_OUT<="0000000000010000";
ELSIF DATA(7 DOWNTO 4) ="1100" THEN
Reg_OUT<="0000000000001000";
ELSIF DATA(7 DOWNTO 4) ="1101" THEN
Reg_OUT<="0000000000000100";
ELSIF DATA(7 DOWNTO 4) ="1110" THEN
Reg_OUT<="0000000000000010";
ELSIF DATA(7 DOWNTO 4) ="1111" THEN
Reg_OUT<="0000000000000001";
END IF;
--
ALU_com<= DATA(15 DOWNTO 12);--THIS VALUE SHOULD EQUAL COMPARE

WHEN BGT3=>   --WAIT
Y_next<= BGT4;
Reg_OUT<=(others =>'0');
ALU_com<=DATA(15 DOWNTO 12);

WHEN BGT4=>

Y_next<=BGT1;
RegG_OUT<='1';

WHEN BGT5=>
y_NEXT<=BGT6;
--Regx_IN
IF DATA(11 DOWNTO 8)="0000" THEN 
Reg_IN<="1000000000000000";
ELSIF DATA(11 DOWNTO 8) ="0001" THEN
Reg_IN<="0100000000000000";
ELSIF DATA(11 DOWNTO 8) ="0010" THEN
Reg_IN<="0010000000000000";
ELSIF DATA(11 DOWNTO 8) ="0011" THEN
Reg_IN<="0001000000000000";
ELSIF DATA(11 DOWNTO 8) ="0100" THEN
Reg_IN<="0000100000000000";
ELSIF DATA(11 DOWNTO 8) ="0101" THEN
Reg_IN<="0000010000000000";
ELSIF DATA(11 DOWNTO 8) ="0110" THEN
Reg_IN<="0000001000000000";
ELSIF DATA(11 DOWNTO 8) ="0111" THEN
Reg_IN<="0000000100000000";
ELSIF DATA(11 DOWNTO 8) ="1000" THEN
Reg_IN<="0000000010000000";
ELSIF DATA(11 DOWNTO 8) ="1001" THEN
Reg_IN<="0000000001000000";
ELSIF DATA(11 DOWNTO 8) ="1010" THEN
Reg_IN<="0000000000100000";
ELSIF DATA(11 DOWNTO 8) ="1011" THEN
Reg_IN<="0000000000010000";
ELSIF DATA(11 DOWNTO 8) ="1100" THEN
Reg_IN<="0000000000001000";
ELSIF DATA(11 DOWNTO 8) ="1101" THEN
Reg_IN<="0000000000000100";
ELSIF DATA(11 DOWNTO 8) ="1110" THEN
Reg_IN<="0000000000000010";
ELSIF DATA(11 DOWNTO 8) ="1111" THEN
Reg_IN<="0000000000000001";
END IF;

WHEN BGT6=>
Y_next<=HOME;
RegG_IN<='0';
RegG_OUT<='0';
Done<='1';




END CASE;
END PROCESS;
END;


